magic
tech sky130A
magscale 1 2
timestamp 1700952384
<< nwell >>
rect 1066 297285 158922 297606
rect 1066 296197 158922 296763
rect 1066 295109 158922 295675
rect 1066 294021 158922 294587
rect 1066 292933 158922 293499
rect 1066 291845 158922 292411
rect 1066 290757 158922 291323
rect 1066 289669 158922 290235
rect 1066 288581 158922 289147
rect 1066 287493 158922 288059
rect 1066 286405 158922 286971
rect 1066 285317 158922 285883
rect 1066 284229 158922 284795
rect 1066 283141 158922 283707
rect 1066 282053 158922 282619
rect 1066 280965 158922 281531
rect 1066 279877 158922 280443
rect 1066 278789 158922 279355
rect 1066 277701 158922 278267
rect 1066 276613 158922 277179
rect 1066 275525 158922 276091
rect 1066 274437 158922 275003
rect 1066 273349 158922 273915
rect 1066 272261 158922 272827
rect 1066 271173 158922 271739
rect 1066 270085 158922 270651
rect 1066 268997 158922 269563
rect 1066 267909 158922 268475
rect 1066 266821 158922 267387
rect 1066 265733 158922 266299
rect 1066 264645 158922 265211
rect 1066 263557 158922 264123
rect 1066 262469 158922 263035
rect 1066 261381 158922 261947
rect 1066 260293 158922 260859
rect 1066 259205 158922 259771
rect 1066 258117 158922 258683
rect 1066 257029 158922 257595
rect 1066 255941 158922 256507
rect 1066 254853 158922 255419
rect 1066 253765 158922 254331
rect 1066 252677 158922 253243
rect 1066 251589 158922 252155
rect 1066 250501 158922 251067
rect 1066 249413 158922 249979
rect 1066 248325 158922 248891
rect 1066 247237 158922 247803
rect 1066 246149 158922 246715
rect 1066 245061 158922 245627
rect 1066 243973 158922 244539
rect 1066 242885 158922 243451
rect 1066 241797 158922 242363
rect 1066 240709 158922 241275
rect 1066 239621 158922 240187
rect 1066 238533 158922 239099
rect 1066 237445 158922 238011
rect 1066 236357 158922 236923
rect 1066 235269 158922 235835
rect 1066 234181 158922 234747
rect 1066 233093 158922 233659
rect 1066 232005 158922 232571
rect 1066 230917 158922 231483
rect 1066 229829 158922 230395
rect 1066 228741 158922 229307
rect 1066 227653 158922 228219
rect 1066 226565 158922 227131
rect 1066 225477 158922 226043
rect 1066 224389 158922 224955
rect 1066 223301 158922 223867
rect 1066 222213 158922 222779
rect 1066 221125 158922 221691
rect 1066 220037 158922 220603
rect 1066 218949 158922 219515
rect 1066 217861 158922 218427
rect 1066 216773 158922 217339
rect 1066 215685 158922 216251
rect 1066 214597 158922 215163
rect 1066 213509 158922 214075
rect 1066 212421 158922 212987
rect 1066 211333 158922 211899
rect 1066 210245 158922 210811
rect 1066 209157 158922 209723
rect 1066 208069 158922 208635
rect 1066 206981 158922 207547
rect 1066 205893 158922 206459
rect 1066 204805 158922 205371
rect 1066 203717 158922 204283
rect 1066 202629 158922 203195
rect 1066 201541 158922 202107
rect 1066 200453 158922 201019
rect 1066 199365 158922 199931
rect 1066 198277 158922 198843
rect 1066 197189 158922 197755
rect 1066 196101 158922 196667
rect 1066 195013 158922 195579
rect 1066 193925 158922 194491
rect 1066 192837 158922 193403
rect 1066 191749 158922 192315
rect 1066 190661 158922 191227
rect 1066 189573 158922 190139
rect 1066 188485 158922 189051
rect 1066 187397 158922 187963
rect 1066 186309 158922 186875
rect 1066 185221 158922 185787
rect 1066 184133 158922 184699
rect 1066 183045 158922 183611
rect 1066 181957 158922 182523
rect 1066 180869 158922 181435
rect 1066 179781 158922 180347
rect 1066 178693 158922 179259
rect 1066 177605 158922 178171
rect 1066 176517 158922 177083
rect 1066 175429 158922 175995
rect 1066 174341 158922 174907
rect 1066 173253 158922 173819
rect 1066 172165 158922 172731
rect 1066 171077 158922 171643
rect 1066 169989 158922 170555
rect 1066 168901 158922 169467
rect 1066 167813 158922 168379
rect 1066 166725 158922 167291
rect 1066 165637 158922 166203
rect 1066 164549 158922 165115
rect 1066 163461 158922 164027
rect 1066 162373 158922 162939
rect 1066 161285 158922 161851
rect 1066 160197 158922 160763
rect 1066 159109 158922 159675
rect 1066 158021 158922 158587
rect 1066 156933 158922 157499
rect 1066 155845 158922 156411
rect 1066 154757 158922 155323
rect 1066 153669 158922 154235
rect 1066 152581 158922 153147
rect 1066 151493 158922 152059
rect 1066 150405 158922 150971
rect 1066 149317 158922 149883
rect 1066 148229 158922 148795
rect 1066 147141 158922 147707
rect 1066 146053 158922 146619
rect 1066 144965 158922 145531
rect 1066 143877 158922 144443
rect 1066 142789 158922 143355
rect 1066 141701 158922 142267
rect 1066 140613 158922 141179
rect 1066 139525 158922 140091
rect 1066 138437 158922 139003
rect 1066 137349 158922 137915
rect 1066 136261 158922 136827
rect 1066 135173 158922 135739
rect 1066 134085 158922 134651
rect 1066 132997 158922 133563
rect 1066 131909 158922 132475
rect 1066 130821 158922 131387
rect 1066 129733 158922 130299
rect 1066 128645 158922 129211
rect 1066 127557 158922 128123
rect 1066 126469 158922 127035
rect 1066 125381 158922 125947
rect 1066 124293 158922 124859
rect 1066 123205 158922 123771
rect 1066 122117 158922 122683
rect 1066 121029 158922 121595
rect 1066 119941 158922 120507
rect 1066 118853 158922 119419
rect 1066 117765 158922 118331
rect 1066 116677 158922 117243
rect 1066 115589 158922 116155
rect 1066 114501 158922 115067
rect 1066 113413 158922 113979
rect 1066 112325 158922 112891
rect 1066 111237 158922 111803
rect 1066 110149 158922 110715
rect 1066 109061 158922 109627
rect 1066 107973 158922 108539
rect 1066 106885 158922 107451
rect 1066 105797 158922 106363
rect 1066 104709 158922 105275
rect 1066 103621 158922 104187
rect 1066 102533 158922 103099
rect 1066 101445 158922 102011
rect 1066 100357 158922 100923
rect 1066 99269 158922 99835
rect 1066 98181 158922 98747
rect 1066 97093 158922 97659
rect 1066 96005 158922 96571
rect 1066 94917 158922 95483
rect 1066 93829 158922 94395
rect 1066 92741 158922 93307
rect 1066 91653 158922 92219
rect 1066 90565 158922 91131
rect 1066 89477 158922 90043
rect 1066 88389 158922 88955
rect 1066 87301 158922 87867
rect 1066 86213 158922 86779
rect 1066 85125 158922 85691
rect 1066 84037 158922 84603
rect 1066 82949 158922 83515
rect 1066 81861 158922 82427
rect 1066 80773 158922 81339
rect 1066 79685 158922 80251
rect 1066 78597 158922 79163
rect 1066 77509 158922 78075
rect 1066 76421 158922 76987
rect 1066 75333 158922 75899
rect 1066 74245 158922 74811
rect 1066 73157 158922 73723
rect 1066 72069 158922 72635
rect 1066 70981 158922 71547
rect 1066 69893 158922 70459
rect 1066 68805 158922 69371
rect 1066 67717 158922 68283
rect 1066 66629 158922 67195
rect 1066 65541 158922 66107
rect 1066 64453 158922 65019
rect 1066 63365 158922 63931
rect 1066 62277 158922 62843
rect 1066 61189 158922 61755
rect 1066 60101 158922 60667
rect 1066 59013 158922 59579
rect 1066 57925 158922 58491
rect 1066 56837 158922 57403
rect 1066 55749 158922 56315
rect 1066 54661 158922 55227
rect 1066 53573 158922 54139
rect 1066 52485 158922 53051
rect 1066 51397 158922 51963
rect 1066 50309 158922 50875
rect 1066 49221 158922 49787
rect 1066 48133 158922 48699
rect 1066 47045 158922 47611
rect 1066 45957 158922 46523
rect 1066 44869 158922 45435
rect 1066 43781 158922 44347
rect 1066 42693 158922 43259
rect 1066 41605 158922 42171
rect 1066 40517 158922 41083
rect 1066 39429 158922 39995
rect 1066 38341 158922 38907
rect 1066 37253 158922 37819
rect 1066 36165 158922 36731
rect 1066 35077 158922 35643
rect 1066 33989 158922 34555
rect 1066 32901 158922 33467
rect 1066 31813 158922 32379
rect 1066 30725 158922 31291
rect 1066 29637 158922 30203
rect 1066 28549 158922 29115
rect 1066 27461 158922 28027
rect 1066 26373 158922 26939
rect 1066 25285 158922 25851
rect 1066 24197 158922 24763
rect 1066 23109 158922 23675
rect 1066 22021 158922 22587
rect 1066 20933 158922 21499
rect 1066 19845 158922 20411
rect 1066 18757 158922 19323
rect 1066 17669 158922 18235
rect 1066 16581 158922 17147
rect 1066 15493 158922 16059
rect 1066 14405 158922 14971
rect 1066 13317 158922 13883
rect 1066 12229 158922 12795
rect 1066 11141 158922 11707
rect 1066 10053 158922 10619
rect 1066 8965 158922 9531
rect 1066 7877 158922 8443
rect 1066 6789 158922 7355
rect 1066 5701 158922 6267
rect 1066 4613 158922 5179
rect 1066 3525 158922 4091
rect 1066 2437 158922 3003
<< obsli1 >>
rect 1104 2159 158884 297585
<< obsm1 >>
rect 1104 2128 158962 297616
<< obsm2 >>
rect 4214 2139 158958 297605
<< metal3 >>
rect 159200 287784 160000 287904
rect 159200 266568 160000 266688
rect 159200 245352 160000 245472
rect 159200 224136 160000 224256
rect 159200 202920 160000 203040
rect 159200 181704 160000 181824
rect 159200 160488 160000 160608
rect 159200 139272 160000 139392
rect 159200 118056 160000 118176
rect 159200 96840 160000 96960
rect 159200 75624 160000 75744
rect 159200 54408 160000 54528
rect 159200 33192 160000 33312
rect 159200 11976 160000 12096
<< obsm3 >>
rect 4210 287984 159200 297601
rect 4210 287704 159120 287984
rect 4210 266768 159200 287704
rect 4210 266488 159120 266768
rect 4210 245552 159200 266488
rect 4210 245272 159120 245552
rect 4210 224336 159200 245272
rect 4210 224056 159120 224336
rect 4210 203120 159200 224056
rect 4210 202840 159120 203120
rect 4210 181904 159200 202840
rect 4210 181624 159120 181904
rect 4210 160688 159200 181624
rect 4210 160408 159120 160688
rect 4210 139472 159200 160408
rect 4210 139192 159120 139472
rect 4210 118256 159200 139192
rect 4210 117976 159120 118256
rect 4210 97040 159200 117976
rect 4210 96760 159120 97040
rect 4210 75824 159200 96760
rect 4210 75544 159120 75824
rect 4210 54608 159200 75544
rect 4210 54328 159120 54608
rect 4210 33392 159200 54328
rect 4210 33112 159120 33392
rect 4210 12176 159200 33112
rect 4210 11896 159120 12176
rect 4210 2143 159200 11896
<< metal4 >>
rect 4208 2128 4528 297616
rect 19568 2128 19888 297616
rect 34928 2128 35248 297616
rect 50288 2128 50608 297616
rect 65648 2128 65968 297616
rect 81008 2128 81328 297616
rect 96368 2128 96688 297616
rect 111728 2128 112048 297616
rect 127088 2128 127408 297616
rect 142448 2128 142768 297616
rect 157808 2128 158128 297616
<< labels >>
rlabel metal3 s 159200 11976 160000 12096 6 clk
port 1 nsew signal input
rlabel metal3 s 159200 160488 160000 160608 6 grant[0]
port 2 nsew signal output
rlabel metal3 s 159200 181704 160000 181824 6 grant[1]
port 3 nsew signal output
rlabel metal3 s 159200 202920 160000 203040 6 grant[2]
port 4 nsew signal output
rlabel metal3 s 159200 224136 160000 224256 6 grant[3]
port 5 nsew signal output
rlabel metal3 s 159200 54408 160000 54528 6 io_oeb[0]
port 6 nsew signal output
rlabel metal3 s 159200 245352 160000 245472 6 io_oeb[1]
port 7 nsew signal output
rlabel metal3 s 159200 266568 160000 266688 6 io_oeb[2]
port 8 nsew signal output
rlabel metal3 s 159200 287784 160000 287904 6 io_oeb[3]
port 9 nsew signal output
rlabel metal3 s 159200 75624 160000 75744 6 req[0]
port 10 nsew signal input
rlabel metal3 s 159200 96840 160000 96960 6 req[1]
port 11 nsew signal input
rlabel metal3 s 159200 118056 160000 118176 6 req[2]
port 12 nsew signal input
rlabel metal3 s 159200 139272 160000 139392 6 req[3]
port 13 nsew signal input
rlabel metal3 s 159200 33192 160000 33312 6 rst
port 14 nsew signal input
rlabel metal4 s 4208 2128 4528 297616 6 vccd1
port 15 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 297616 6 vccd1
port 15 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 297616 6 vccd1
port 15 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 297616 6 vccd1
port 15 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 297616 6 vccd1
port 15 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 297616 6 vccd1
port 15 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 297616 6 vssd1
port 16 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 297616 6 vssd1
port 16 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 297616 6 vssd1
port 16 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 297616 6 vssd1
port 16 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 297616 6 vssd1
port 16 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 160000 300000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 12816210
string GDS_FILE /home/navya/asic_project/pes_rr_arbiter_tapeout/openlane/pes_rr_arbiter/runs/23_11_26_04_12/results/signoff/pes_rr_arbiter.magic.gds
string GDS_START 215348
<< end >>

