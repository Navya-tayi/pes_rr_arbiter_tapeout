VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO pes_rr_arbiter
  CLASS BLOCK ;
  FOREIGN pes_rr_arbiter ;
  ORIGIN 0.000 0.000 ;
  SIZE 800.000 BY 1500.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 796.000 59.880 800.000 60.480 ;
    END
  END clk
  PIN grant[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 802.440 800.000 803.040 ;
    END
  END grant[0]
  PIN grant[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 908.520 800.000 909.120 ;
    END
  END grant[1]
  PIN grant[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1014.600 800.000 1015.200 ;
    END
  END grant[2]
  PIN grant[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1120.680 800.000 1121.280 ;
    END
  END grant[3]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 272.040 800.000 272.640 ;
    END
  END io_oeb[0]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1226.760 800.000 1227.360 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1332.840 800.000 1333.440 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 1438.920 800.000 1439.520 ;
    END
  END io_oeb[3]
  PIN req[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 378.120 800.000 378.720 ;
    END
  END req[0]
  PIN req[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 484.200 800.000 484.800 ;
    END
  END req[1]
  PIN req[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 590.280 800.000 590.880 ;
    END
  END req[2]
  PIN req[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 696.360 800.000 696.960 ;
    END
  END req[3]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 165.960 800.000 166.560 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1488.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1488.080 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 1486.425 794.610 1488.030 ;
        RECT 5.330 1480.985 794.610 1483.815 ;
        RECT 5.330 1475.545 794.610 1478.375 ;
        RECT 5.330 1470.105 794.610 1472.935 ;
        RECT 5.330 1464.665 794.610 1467.495 ;
        RECT 5.330 1459.225 794.610 1462.055 ;
        RECT 5.330 1453.785 794.610 1456.615 ;
        RECT 5.330 1448.345 794.610 1451.175 ;
        RECT 5.330 1442.905 794.610 1445.735 ;
        RECT 5.330 1437.465 794.610 1440.295 ;
        RECT 5.330 1432.025 794.610 1434.855 ;
        RECT 5.330 1426.585 794.610 1429.415 ;
        RECT 5.330 1421.145 794.610 1423.975 ;
        RECT 5.330 1415.705 794.610 1418.535 ;
        RECT 5.330 1410.265 794.610 1413.095 ;
        RECT 5.330 1404.825 794.610 1407.655 ;
        RECT 5.330 1399.385 794.610 1402.215 ;
        RECT 5.330 1393.945 794.610 1396.775 ;
        RECT 5.330 1388.505 794.610 1391.335 ;
        RECT 5.330 1383.065 794.610 1385.895 ;
        RECT 5.330 1377.625 794.610 1380.455 ;
        RECT 5.330 1372.185 794.610 1375.015 ;
        RECT 5.330 1366.745 794.610 1369.575 ;
        RECT 5.330 1361.305 794.610 1364.135 ;
        RECT 5.330 1355.865 794.610 1358.695 ;
        RECT 5.330 1350.425 794.610 1353.255 ;
        RECT 5.330 1344.985 794.610 1347.815 ;
        RECT 5.330 1339.545 794.610 1342.375 ;
        RECT 5.330 1334.105 794.610 1336.935 ;
        RECT 5.330 1328.665 794.610 1331.495 ;
        RECT 5.330 1323.225 794.610 1326.055 ;
        RECT 5.330 1317.785 794.610 1320.615 ;
        RECT 5.330 1312.345 794.610 1315.175 ;
        RECT 5.330 1306.905 794.610 1309.735 ;
        RECT 5.330 1301.465 794.610 1304.295 ;
        RECT 5.330 1296.025 794.610 1298.855 ;
        RECT 5.330 1290.585 794.610 1293.415 ;
        RECT 5.330 1285.145 794.610 1287.975 ;
        RECT 5.330 1279.705 794.610 1282.535 ;
        RECT 5.330 1274.265 794.610 1277.095 ;
        RECT 5.330 1268.825 794.610 1271.655 ;
        RECT 5.330 1263.385 794.610 1266.215 ;
        RECT 5.330 1257.945 794.610 1260.775 ;
        RECT 5.330 1252.505 794.610 1255.335 ;
        RECT 5.330 1247.065 794.610 1249.895 ;
        RECT 5.330 1241.625 794.610 1244.455 ;
        RECT 5.330 1236.185 794.610 1239.015 ;
        RECT 5.330 1230.745 794.610 1233.575 ;
        RECT 5.330 1225.305 794.610 1228.135 ;
        RECT 5.330 1219.865 794.610 1222.695 ;
        RECT 5.330 1214.425 794.610 1217.255 ;
        RECT 5.330 1208.985 794.610 1211.815 ;
        RECT 5.330 1203.545 794.610 1206.375 ;
        RECT 5.330 1198.105 794.610 1200.935 ;
        RECT 5.330 1192.665 794.610 1195.495 ;
        RECT 5.330 1187.225 794.610 1190.055 ;
        RECT 5.330 1181.785 794.610 1184.615 ;
        RECT 5.330 1176.345 794.610 1179.175 ;
        RECT 5.330 1170.905 794.610 1173.735 ;
        RECT 5.330 1165.465 794.610 1168.295 ;
        RECT 5.330 1160.025 794.610 1162.855 ;
        RECT 5.330 1154.585 794.610 1157.415 ;
        RECT 5.330 1149.145 794.610 1151.975 ;
        RECT 5.330 1143.705 794.610 1146.535 ;
        RECT 5.330 1138.265 794.610 1141.095 ;
        RECT 5.330 1132.825 794.610 1135.655 ;
        RECT 5.330 1127.385 794.610 1130.215 ;
        RECT 5.330 1121.945 794.610 1124.775 ;
        RECT 5.330 1116.505 794.610 1119.335 ;
        RECT 5.330 1111.065 794.610 1113.895 ;
        RECT 5.330 1105.625 794.610 1108.455 ;
        RECT 5.330 1100.185 794.610 1103.015 ;
        RECT 5.330 1094.745 794.610 1097.575 ;
        RECT 5.330 1089.305 794.610 1092.135 ;
        RECT 5.330 1083.865 794.610 1086.695 ;
        RECT 5.330 1078.425 794.610 1081.255 ;
        RECT 5.330 1072.985 794.610 1075.815 ;
        RECT 5.330 1067.545 794.610 1070.375 ;
        RECT 5.330 1062.105 794.610 1064.935 ;
        RECT 5.330 1056.665 794.610 1059.495 ;
        RECT 5.330 1051.225 794.610 1054.055 ;
        RECT 5.330 1045.785 794.610 1048.615 ;
        RECT 5.330 1040.345 794.610 1043.175 ;
        RECT 5.330 1034.905 794.610 1037.735 ;
        RECT 5.330 1029.465 794.610 1032.295 ;
        RECT 5.330 1024.025 794.610 1026.855 ;
        RECT 5.330 1018.585 794.610 1021.415 ;
        RECT 5.330 1013.145 794.610 1015.975 ;
        RECT 5.330 1007.705 794.610 1010.535 ;
        RECT 5.330 1002.265 794.610 1005.095 ;
        RECT 5.330 996.825 794.610 999.655 ;
        RECT 5.330 991.385 794.610 994.215 ;
        RECT 5.330 985.945 794.610 988.775 ;
        RECT 5.330 980.505 794.610 983.335 ;
        RECT 5.330 975.065 794.610 977.895 ;
        RECT 5.330 969.625 794.610 972.455 ;
        RECT 5.330 964.185 794.610 967.015 ;
        RECT 5.330 958.745 794.610 961.575 ;
        RECT 5.330 953.305 794.610 956.135 ;
        RECT 5.330 947.865 794.610 950.695 ;
        RECT 5.330 942.425 794.610 945.255 ;
        RECT 5.330 936.985 794.610 939.815 ;
        RECT 5.330 931.545 794.610 934.375 ;
        RECT 5.330 926.105 794.610 928.935 ;
        RECT 5.330 920.665 794.610 923.495 ;
        RECT 5.330 915.225 794.610 918.055 ;
        RECT 5.330 909.785 794.610 912.615 ;
        RECT 5.330 904.345 794.610 907.175 ;
        RECT 5.330 898.905 794.610 901.735 ;
        RECT 5.330 893.465 794.610 896.295 ;
        RECT 5.330 888.025 794.610 890.855 ;
        RECT 5.330 882.585 794.610 885.415 ;
        RECT 5.330 877.145 794.610 879.975 ;
        RECT 5.330 871.705 794.610 874.535 ;
        RECT 5.330 866.265 794.610 869.095 ;
        RECT 5.330 860.825 794.610 863.655 ;
        RECT 5.330 855.385 794.610 858.215 ;
        RECT 5.330 849.945 794.610 852.775 ;
        RECT 5.330 844.505 794.610 847.335 ;
        RECT 5.330 839.065 794.610 841.895 ;
        RECT 5.330 833.625 794.610 836.455 ;
        RECT 5.330 828.185 794.610 831.015 ;
        RECT 5.330 822.745 794.610 825.575 ;
        RECT 5.330 817.305 794.610 820.135 ;
        RECT 5.330 811.865 794.610 814.695 ;
        RECT 5.330 806.425 794.610 809.255 ;
        RECT 5.330 800.985 794.610 803.815 ;
        RECT 5.330 795.545 794.610 798.375 ;
        RECT 5.330 790.105 794.610 792.935 ;
        RECT 5.330 784.665 794.610 787.495 ;
        RECT 5.330 779.225 794.610 782.055 ;
        RECT 5.330 773.785 794.610 776.615 ;
        RECT 5.330 768.345 794.610 771.175 ;
        RECT 5.330 762.905 794.610 765.735 ;
        RECT 5.330 757.465 794.610 760.295 ;
        RECT 5.330 752.025 794.610 754.855 ;
        RECT 5.330 746.585 794.610 749.415 ;
        RECT 5.330 741.145 794.610 743.975 ;
        RECT 5.330 735.705 794.610 738.535 ;
        RECT 5.330 730.265 794.610 733.095 ;
        RECT 5.330 724.825 794.610 727.655 ;
        RECT 5.330 719.385 794.610 722.215 ;
        RECT 5.330 713.945 794.610 716.775 ;
        RECT 5.330 708.505 794.610 711.335 ;
        RECT 5.330 703.065 794.610 705.895 ;
        RECT 5.330 697.625 794.610 700.455 ;
        RECT 5.330 692.185 794.610 695.015 ;
        RECT 5.330 686.745 794.610 689.575 ;
        RECT 5.330 681.305 794.610 684.135 ;
        RECT 5.330 675.865 794.610 678.695 ;
        RECT 5.330 670.425 794.610 673.255 ;
        RECT 5.330 664.985 794.610 667.815 ;
        RECT 5.330 659.545 794.610 662.375 ;
        RECT 5.330 654.105 794.610 656.935 ;
        RECT 5.330 648.665 794.610 651.495 ;
        RECT 5.330 643.225 794.610 646.055 ;
        RECT 5.330 637.785 794.610 640.615 ;
        RECT 5.330 632.345 794.610 635.175 ;
        RECT 5.330 626.905 794.610 629.735 ;
        RECT 5.330 621.465 794.610 624.295 ;
        RECT 5.330 616.025 794.610 618.855 ;
        RECT 5.330 610.585 794.610 613.415 ;
        RECT 5.330 605.145 794.610 607.975 ;
        RECT 5.330 599.705 794.610 602.535 ;
        RECT 5.330 594.265 794.610 597.095 ;
        RECT 5.330 588.825 794.610 591.655 ;
        RECT 5.330 583.385 794.610 586.215 ;
        RECT 5.330 577.945 794.610 580.775 ;
        RECT 5.330 572.505 794.610 575.335 ;
        RECT 5.330 567.065 794.610 569.895 ;
        RECT 5.330 561.625 794.610 564.455 ;
        RECT 5.330 556.185 794.610 559.015 ;
        RECT 5.330 550.745 794.610 553.575 ;
        RECT 5.330 545.305 794.610 548.135 ;
        RECT 5.330 539.865 794.610 542.695 ;
        RECT 5.330 534.425 794.610 537.255 ;
        RECT 5.330 528.985 794.610 531.815 ;
        RECT 5.330 523.545 794.610 526.375 ;
        RECT 5.330 518.105 794.610 520.935 ;
        RECT 5.330 512.665 794.610 515.495 ;
        RECT 5.330 507.225 794.610 510.055 ;
        RECT 5.330 501.785 794.610 504.615 ;
        RECT 5.330 496.345 794.610 499.175 ;
        RECT 5.330 490.905 794.610 493.735 ;
        RECT 5.330 485.465 794.610 488.295 ;
        RECT 5.330 480.025 794.610 482.855 ;
        RECT 5.330 474.585 794.610 477.415 ;
        RECT 5.330 469.145 794.610 471.975 ;
        RECT 5.330 463.705 794.610 466.535 ;
        RECT 5.330 458.265 794.610 461.095 ;
        RECT 5.330 452.825 794.610 455.655 ;
        RECT 5.330 447.385 794.610 450.215 ;
        RECT 5.330 441.945 794.610 444.775 ;
        RECT 5.330 436.505 794.610 439.335 ;
        RECT 5.330 431.065 794.610 433.895 ;
        RECT 5.330 425.625 794.610 428.455 ;
        RECT 5.330 420.185 794.610 423.015 ;
        RECT 5.330 414.745 794.610 417.575 ;
        RECT 5.330 409.305 794.610 412.135 ;
        RECT 5.330 403.865 794.610 406.695 ;
        RECT 5.330 398.425 794.610 401.255 ;
        RECT 5.330 392.985 794.610 395.815 ;
        RECT 5.330 387.545 794.610 390.375 ;
        RECT 5.330 382.105 794.610 384.935 ;
        RECT 5.330 376.665 794.610 379.495 ;
        RECT 5.330 371.225 794.610 374.055 ;
        RECT 5.330 365.785 794.610 368.615 ;
        RECT 5.330 360.345 794.610 363.175 ;
        RECT 5.330 354.905 794.610 357.735 ;
        RECT 5.330 349.465 794.610 352.295 ;
        RECT 5.330 344.025 794.610 346.855 ;
        RECT 5.330 338.585 794.610 341.415 ;
        RECT 5.330 333.145 794.610 335.975 ;
        RECT 5.330 327.705 794.610 330.535 ;
        RECT 5.330 322.265 794.610 325.095 ;
        RECT 5.330 316.825 794.610 319.655 ;
        RECT 5.330 311.385 794.610 314.215 ;
        RECT 5.330 305.945 794.610 308.775 ;
        RECT 5.330 300.505 794.610 303.335 ;
        RECT 5.330 295.065 794.610 297.895 ;
        RECT 5.330 289.625 794.610 292.455 ;
        RECT 5.330 284.185 794.610 287.015 ;
        RECT 5.330 278.745 794.610 281.575 ;
        RECT 5.330 273.305 794.610 276.135 ;
        RECT 5.330 267.865 794.610 270.695 ;
        RECT 5.330 262.425 794.610 265.255 ;
        RECT 5.330 256.985 794.610 259.815 ;
        RECT 5.330 251.545 794.610 254.375 ;
        RECT 5.330 246.105 794.610 248.935 ;
        RECT 5.330 240.665 794.610 243.495 ;
        RECT 5.330 235.225 794.610 238.055 ;
        RECT 5.330 229.785 794.610 232.615 ;
        RECT 5.330 224.345 794.610 227.175 ;
        RECT 5.330 218.905 794.610 221.735 ;
        RECT 5.330 213.465 794.610 216.295 ;
        RECT 5.330 208.025 794.610 210.855 ;
        RECT 5.330 202.585 794.610 205.415 ;
        RECT 5.330 197.145 794.610 199.975 ;
        RECT 5.330 191.705 794.610 194.535 ;
        RECT 5.330 186.265 794.610 189.095 ;
        RECT 5.330 180.825 794.610 183.655 ;
        RECT 5.330 175.385 794.610 178.215 ;
        RECT 5.330 169.945 794.610 172.775 ;
        RECT 5.330 164.505 794.610 167.335 ;
        RECT 5.330 159.065 794.610 161.895 ;
        RECT 5.330 153.625 794.610 156.455 ;
        RECT 5.330 148.185 794.610 151.015 ;
        RECT 5.330 142.745 794.610 145.575 ;
        RECT 5.330 137.305 794.610 140.135 ;
        RECT 5.330 131.865 794.610 134.695 ;
        RECT 5.330 126.425 794.610 129.255 ;
        RECT 5.330 120.985 794.610 123.815 ;
        RECT 5.330 115.545 794.610 118.375 ;
        RECT 5.330 110.105 794.610 112.935 ;
        RECT 5.330 104.665 794.610 107.495 ;
        RECT 5.330 99.225 794.610 102.055 ;
        RECT 5.330 93.785 794.610 96.615 ;
        RECT 5.330 88.345 794.610 91.175 ;
        RECT 5.330 82.905 794.610 85.735 ;
        RECT 5.330 77.465 794.610 80.295 ;
        RECT 5.330 72.025 794.610 74.855 ;
        RECT 5.330 66.585 794.610 69.415 ;
        RECT 5.330 61.145 794.610 63.975 ;
        RECT 5.330 55.705 794.610 58.535 ;
        RECT 5.330 50.265 794.610 53.095 ;
        RECT 5.330 44.825 794.610 47.655 ;
        RECT 5.330 39.385 794.610 42.215 ;
        RECT 5.330 33.945 794.610 36.775 ;
        RECT 5.330 28.505 794.610 31.335 ;
        RECT 5.330 23.065 794.610 25.895 ;
        RECT 5.330 17.625 794.610 20.455 ;
        RECT 5.330 12.185 794.610 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 794.420 1487.925 ;
      LAYER met1 ;
        RECT 5.520 10.640 794.810 1488.080 ;
      LAYER met2 ;
        RECT 21.070 10.695 794.790 1488.025 ;
      LAYER met3 ;
        RECT 21.050 1439.920 796.000 1488.005 ;
        RECT 21.050 1438.520 795.600 1439.920 ;
        RECT 21.050 1333.840 796.000 1438.520 ;
        RECT 21.050 1332.440 795.600 1333.840 ;
        RECT 21.050 1227.760 796.000 1332.440 ;
        RECT 21.050 1226.360 795.600 1227.760 ;
        RECT 21.050 1121.680 796.000 1226.360 ;
        RECT 21.050 1120.280 795.600 1121.680 ;
        RECT 21.050 1015.600 796.000 1120.280 ;
        RECT 21.050 1014.200 795.600 1015.600 ;
        RECT 21.050 909.520 796.000 1014.200 ;
        RECT 21.050 908.120 795.600 909.520 ;
        RECT 21.050 803.440 796.000 908.120 ;
        RECT 21.050 802.040 795.600 803.440 ;
        RECT 21.050 697.360 796.000 802.040 ;
        RECT 21.050 695.960 795.600 697.360 ;
        RECT 21.050 591.280 796.000 695.960 ;
        RECT 21.050 589.880 795.600 591.280 ;
        RECT 21.050 485.200 796.000 589.880 ;
        RECT 21.050 483.800 795.600 485.200 ;
        RECT 21.050 379.120 796.000 483.800 ;
        RECT 21.050 377.720 795.600 379.120 ;
        RECT 21.050 273.040 796.000 377.720 ;
        RECT 21.050 271.640 795.600 273.040 ;
        RECT 21.050 166.960 796.000 271.640 ;
        RECT 21.050 165.560 795.600 166.960 ;
        RECT 21.050 60.880 796.000 165.560 ;
        RECT 21.050 59.480 795.600 60.880 ;
        RECT 21.050 10.715 796.000 59.480 ;
  END
END pes_rr_arbiter
END LIBRARY

